// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none

`timescale 1 ns / 1 ps

`include "udp_host.v"
`include "uprj_netlists.v"
`include "caravel_netlists.v"
`include "spiflash.v"

module ethernet_100m_tb;
	reg clock;
	reg RSTB;
	reg CSB;
	reg power1, power2;
	reg power3, power4;

	wire gpio;
	wire [37:0] mprj_io;
	
	reg  rst;
	wire [3:0] phy_txd;
    wire phy_tx_en;
    wire phy_tx_clk;
    wire phy_rx_clk;
    wire [3:0] phy_rxd;
    wire phy_rx_dv;
    wire phy_rx_er;

    integer clock_counter = 0;
    integer f = 0;

    assign mprj_io[8]	= rst;
	assign phy_txd		= mprj_io[21:18];
    assign phy_tx_en	= mprj_io[17];
    assign phy_tx_clk	= mprj_io[16];
    assign phy_rx_clk	= mprj_io[9];
    assign phy_rxd 		= mprj_io[15:12];
    assign phy_rx_dv	= mprj_io[10];
    assign phy_rx_er	= mprj_io[11];

	assign mprj_io[3] = (CSB == 1'b1) ? 1'b1 : 1'bz;

	// External clock is used by default.  Make this artificially fast for the
	// simulation.  Normally this would be a slow clock and the digital PLL
	// would be the fast clock.

	always #20 clock <= (clock === 1'b0);

	always @(posedge clock) begin
		clock_counter = clock_counter + 1;
		if (clock_counter == 25) $fwrite(f, "%d nanoseconds elapsed.\n", clock_counter*40);
	end

	initial begin
	   clock = 0;
	   rst = 0;

	   f = $fopen("output.txt","w");
	   $fwrite(f, "Test Ethernet 100Mbps Started");

	   #172001 wait(CSB);
	   
	   #1000 rst = 1;
	   #100  rst = 0;

	   #100000;
	   `ifdef GL
	      $display ("Monitor: Timeout, Test Ethernet 100Mbps (GL) Failed");
	   `else
	      $display ("Monitor: Timeout, Test Ethernet 100Mbps (RTL) Failed");
	   `endif
	   $finish;
	end

	initial begin
		RSTB <= 1'b0;
		CSB  <= 1'b1;		// Force CSB high
		#2000;
		RSTB <= 1'b1;	    	// Release reset
		#170000;
		CSB = 1'b0;		// CSB can be released
	end

	initial begin		// Power-up sequence
		power1 <= 1'b0;
		power2 <= 1'b0;
		power3 <= 1'b0;
		power4 <= 1'b0;
		#100;
		power1 <= 1'b1;
		#100;
		power2 <= 1'b1;
		#100;
		power3 <= 1'b1;
		#100;
		power4 <= 1'b1;
	end

	always @(mprj_io) begin
		#1 $display("MPRJ-IO state = %b ", mprj_io[7:0]);
	end

	wire flash_csb;
	wire flash_clk;
	wire flash_io0;
	wire flash_io1;

	wire VDD3V3 = power1;
	wire VDD1V8 = power2;
	wire USER_VDD3V3 = power3;
	wire USER_VDD1V8 = power4;
	wire VSS = 1'b0;

	udp_host host(
	    .clk(clock),
	    .rst(rst),
	    .phy_txd(phy_txd),
	    .phy_tx_en(phy_tx_en),
	    .phy_tx_clk(phy_tx_clk),
	    .phy_rx_clk(phy_rx_clk),
	    .phy_rxd(phy_rxd),
	    .phy_rx_dv(phy_rx_dv),
	    .phy_rx_er(phy_rx_er)
    );

	caravel uut (
		.vddio	  (VDD3V3),
		.vssio	  (VSS),
		.vdda	  (VDD3V3),
		.vssa	  (VSS),
		.vccd	  (VDD1V8),
		.vssd	  (VSS),
		.vdda1    (USER_VDD3V3),
		.vdda2    (USER_VDD3V3),
		.vssa1	  (VSS),
		.vssa2	  (VSS),
		.vccd1	  (USER_VDD1V8),
		.vccd2	  (USER_VDD1V8),
		.vssd1	  (VSS),
		.vssd2	  (VSS),
		.clock	  (clock),
		.gpio     (gpio),
        .mprj_io  (mprj_io),
		.flash_csb(flash_csb),
		.flash_clk(flash_clk),
		.flash_io0(flash_io0),
		.flash_io1(flash_io1),
		.resetb	  (RSTB)
	);

	spiflash #(
		.FILENAME("ethernet_100m.hex")
	) spiflash (
		.csb(flash_csb),
		.clk(flash_clk),
		.io0(flash_io0),
		.io1(flash_io1),
		.io2(),			// not used
		.io3()			// not used
	);

endmodule
`default_nettype wire